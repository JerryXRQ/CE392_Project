// RFS_WiFi.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module RFS_WiFi (
		input  wire        clk_clk,                                   //                                clk.clk
		input  wire [11:0] pio_height_external_connection_export,     //     pio_height_external_connection.export
		input  wire [1:0]  pio_key_external_connection_export,        //        pio_key_external_connection.export
		output wire [3:0]  pio_led_external_connection_export,        //        pio_led_external_connection.export
		input  wire [11:0] pio_width_external_connection_export,      //      pio_width_external_connection.export
		output wire        pio_wifi_reset_external_connection_export, // pio_wifi_reset_external_connection.export
		input  wire [11:0] pio_x_external_connection_export,          //          pio_x_external_connection.export
		input  wire [11:0] pio_y_external_connection_export,          //          pio_y_external_connection.export
		input  wire        reset_reset_n,                             //                              reset.reset_n
		output wire [47:0] seg7_if_0_conduit_end_export,              //              seg7_if_0_conduit_end.export
		input  wire        wifi_uart0_external_connection_rxd,        //     wifi_uart0_external_connection.rxd
		output wire        wifi_uart0_external_connection_txd,        //                                   .txd
		input  wire        wifi_uart0_external_connection_cts_n,      //                                   .cts_n
		output wire        wifi_uart0_external_connection_rts_n       //                                   .rts_n
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                          // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                       // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                       // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [19:0] nios2_gen2_0_data_master_address;                           // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                        // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                              // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                     // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                             // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                         // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                   // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [19:0] nios2_gen2_0_instruction_master_address;                    // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                       // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;              // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;     // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;  // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [7:0] mm_interconnect_0_seg7_if_0_avalon_slave_readdata;          // SEG7_IF_0:s_readdata -> mm_interconnect_0:SEG7_IF_0_avalon_slave_readdata
	wire   [2:0] mm_interconnect_0_seg7_if_0_avalon_slave_address;           // mm_interconnect_0:SEG7_IF_0_avalon_slave_address -> SEG7_IF_0:s_address
	wire         mm_interconnect_0_seg7_if_0_avalon_slave_read;              // mm_interconnect_0:SEG7_IF_0_avalon_slave_read -> SEG7_IF_0:s_read
	wire         mm_interconnect_0_seg7_if_0_avalon_slave_write;             // mm_interconnect_0:SEG7_IF_0_avalon_slave_write -> SEG7_IF_0:s_write
	wire   [7:0] mm_interconnect_0_seg7_if_0_avalon_slave_writedata;         // mm_interconnect_0:SEG7_IF_0_avalon_slave_writedata -> SEG7_IF_0:s_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;        // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;         // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;    // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest; // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_timer_s1_chipselect;                      // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                        // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                         // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                           // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                       // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_pio_key_s1_chipselect;                    // mm_interconnect_0:pio_key_s1_chipselect -> pio_key:chipselect
	wire  [31:0] mm_interconnect_0_pio_key_s1_readdata;                      // pio_key:readdata -> mm_interconnect_0:pio_key_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_key_s1_address;                       // mm_interconnect_0:pio_key_s1_address -> pio_key:address
	wire         mm_interconnect_0_pio_key_s1_write;                         // mm_interconnect_0:pio_key_s1_write -> pio_key:write_n
	wire  [31:0] mm_interconnect_0_pio_key_s1_writedata;                     // mm_interconnect_0:pio_key_s1_writedata -> pio_key:writedata
	wire         mm_interconnect_0_wifi_uart0_s1_chipselect;                 // mm_interconnect_0:wifi_uart0_s1_chipselect -> wifi_uart0:chipselect
	wire  [15:0] mm_interconnect_0_wifi_uart0_s1_readdata;                   // wifi_uart0:readdata -> mm_interconnect_0:wifi_uart0_s1_readdata
	wire   [2:0] mm_interconnect_0_wifi_uart0_s1_address;                    // mm_interconnect_0:wifi_uart0_s1_address -> wifi_uart0:address
	wire         mm_interconnect_0_wifi_uart0_s1_read;                       // mm_interconnect_0:wifi_uart0_s1_read -> wifi_uart0:read_n
	wire         mm_interconnect_0_wifi_uart0_s1_begintransfer;              // mm_interconnect_0:wifi_uart0_s1_begintransfer -> wifi_uart0:begintransfer
	wire         mm_interconnect_0_wifi_uart0_s1_write;                      // mm_interconnect_0:wifi_uart0_s1_write -> wifi_uart0:write_n
	wire  [15:0] mm_interconnect_0_wifi_uart0_s1_writedata;                  // mm_interconnect_0:wifi_uart0_s1_writedata -> wifi_uart0:writedata
	wire         mm_interconnect_0_pio_wifi_reset_s1_chipselect;             // mm_interconnect_0:pio_wifi_reset_s1_chipselect -> pio_wifi_reset:chipselect
	wire  [31:0] mm_interconnect_0_pio_wifi_reset_s1_readdata;               // pio_wifi_reset:readdata -> mm_interconnect_0:pio_wifi_reset_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_wifi_reset_s1_address;                // mm_interconnect_0:pio_wifi_reset_s1_address -> pio_wifi_reset:address
	wire         mm_interconnect_0_pio_wifi_reset_s1_write;                  // mm_interconnect_0:pio_wifi_reset_s1_write -> pio_wifi_reset:write_n
	wire  [31:0] mm_interconnect_0_pio_wifi_reset_s1_writedata;              // mm_interconnect_0:pio_wifi_reset_s1_writedata -> pio_wifi_reset:writedata
	wire         mm_interconnect_0_pio_led_s1_chipselect;                    // mm_interconnect_0:pio_led_s1_chipselect -> pio_led:chipselect
	wire  [31:0] mm_interconnect_0_pio_led_s1_readdata;                      // pio_led:readdata -> mm_interconnect_0:pio_led_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_led_s1_address;                       // mm_interconnect_0:pio_led_s1_address -> pio_led:address
	wire         mm_interconnect_0_pio_led_s1_write;                         // mm_interconnect_0:pio_led_s1_write -> pio_led:write_n
	wire  [31:0] mm_interconnect_0_pio_led_s1_writedata;                     // mm_interconnect_0:pio_led_s1_writedata -> pio_led:writedata
	wire  [31:0] mm_interconnect_0_pio_x_s1_readdata;                        // pio_x:readdata -> mm_interconnect_0:pio_x_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_x_s1_address;                         // mm_interconnect_0:pio_x_s1_address -> pio_x:address
	wire  [31:0] mm_interconnect_0_pio_y_s1_readdata;                        // pio_y:readdata -> mm_interconnect_0:pio_y_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_y_s1_address;                         // mm_interconnect_0:pio_y_s1_address -> pio_y:address
	wire  [31:0] mm_interconnect_0_pio_width_s1_readdata;                    // pio_width:readdata -> mm_interconnect_0:pio_width_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_width_s1_address;                     // mm_interconnect_0:pio_width_s1_address -> pio_width:address
	wire  [31:0] mm_interconnect_0_pio_height_s1_readdata;                   // pio_height:readdata -> mm_interconnect_0:pio_height_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_height_s1_address;                    // mm_interconnect_0:pio_height_s1_address -> pio_height:address
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;             // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;               // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_s1_address;                // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;             // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                  // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;              // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                  // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         irq_mapper_receiver0_irq;                                   // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                   // timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                   // pio_key:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                   // wifi_uart0:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                       // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [SEG7_IF_0:s_reset, jtag_uart:rst_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, onchip_memory2:reset, pio_height:reset_n, pio_key:reset_n, pio_led:reset_n, pio_width:reset_n, pio_wifi_reset:reset_n, pio_x:reset_n, pio_y:reset_n, rst_translator:in_reset, sysid_qsys:reset_n, timer:reset_n, wifi_uart0:reset_n]
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [onchip_memory2:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                     // rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, rst_translator_001:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                     // nios2_gen2_0:debug_reset_request -> rst_controller_001:reset_in1

	SEG7_IF #(
		.SEG7_NUM       (6),
		.ADDR_WIDTH     (3),
		.DEFAULT_ACTIVE (1),
		.LOW_ACTIVE     (1)
	) seg7_if_0 (
		.s_address   (mm_interconnect_0_seg7_if_0_avalon_slave_address),   //     avalon_slave.address
		.s_read      (mm_interconnect_0_seg7_if_0_avalon_slave_read),      //                 .read
		.s_readdata  (mm_interconnect_0_seg7_if_0_avalon_slave_readdata),  //                 .readdata
		.s_write     (mm_interconnect_0_seg7_if_0_avalon_slave_write),     //                 .write
		.s_writedata (mm_interconnect_0_seg7_if_0_avalon_slave_writedata), //                 .writedata
		.SEG7        (seg7_if_0_conduit_end_export),                       //      conduit_end.export
		.s_clk       (clk_clk),                                            //       clock_sink.clk
		.s_reset     (rst_controller_reset_out_reset)                      // clock_sink_reset.reset
	);

	RFS_WiFi_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	RFS_WiFi_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	RFS_WiFi_onchip_memory2 onchip_memory2 (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	RFS_WiFi_pio_height pio_height (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_pio_height_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_height_s1_readdata), //                    .readdata
		.in_port  (pio_height_external_connection_export)     // external_connection.export
	);

	RFS_WiFi_pio_key pio_key (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_key_s1_readdata),   //                    .readdata
		.in_port    (pio_key_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                 //                 irq.irq
	);

	RFS_WiFi_pio_led pio_led (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_s1_readdata),   //                    .readdata
		.out_port   (pio_led_external_connection_export)       // external_connection.export
	);

	RFS_WiFi_pio_height pio_width (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_pio_width_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_width_s1_readdata), //                    .readdata
		.in_port  (pio_width_external_connection_export)     // external_connection.export
	);

	RFS_WiFi_pio_wifi_reset pio_wifi_reset (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_pio_wifi_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_wifi_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_wifi_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_wifi_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_wifi_reset_s1_readdata),   //                    .readdata
		.out_port   (pio_wifi_reset_external_connection_export)       // external_connection.export
	);

	RFS_WiFi_pio_height pio_x (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_pio_x_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_x_s1_readdata), //                    .readdata
		.in_port  (pio_x_external_connection_export)     // external_connection.export
	);

	RFS_WiFi_pio_height pio_y (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_pio_y_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_y_s1_readdata), //                    .readdata
		.in_port  (pio_y_external_connection_export)     // external_connection.export
	);

	RFS_WiFi_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	RFS_WiFi_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	RFS_WiFi_wifi_uart0 wifi_uart0 (
		.clk           (clk_clk),                                       //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address       (mm_interconnect_0_wifi_uart0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_wifi_uart0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_wifi_uart0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_wifi_uart0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_wifi_uart0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_wifi_uart0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_wifi_uart0_s1_readdata),      //                    .readdata
		.rxd           (wifi_uart0_external_connection_rxd),            // external_connection.export
		.txd           (wifi_uart0_external_connection_txd),            //                    .export
		.cts_n         (wifi_uart0_external_connection_cts_n),          //                    .export
		.rts_n         (wifi_uart0_external_connection_rts_n),          //                    .export
		.irq           (irq_mapper_receiver3_irq)                       //                 irq.irq
	);

	RFS_WiFi_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                 (clk_clk),                                                    //                               clk_50_clk.clk
		.jtag_uart_reset_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                             //    jtag_uart_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                         // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                           //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                       //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                        //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                              //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                          //                                         .readdata
		.nios2_gen2_0_data_master_readdatavalid         (nios2_gen2_0_data_master_readdatavalid),                     //                                         .readdatavalid
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                             //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                         //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                       //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                    //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                       //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                   //                                         .readdata
		.nios2_gen2_0_instruction_master_readdatavalid  (nios2_gen2_0_instruction_master_readdatavalid),              //                                         .readdatavalid
		.jtag_uart_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),      //              jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),        //                                         .write
		.jtag_uart_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),         //                                         .read
		.jtag_uart_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),     //                                         .readdata
		.jtag_uart_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),    //                                         .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),  //                                         .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),   //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                                         .debugaccess
		.onchip_memory2_s1_address                      (mm_interconnect_0_onchip_memory2_s1_address),                //                        onchip_memory2_s1.address
		.onchip_memory2_s1_write                        (mm_interconnect_0_onchip_memory2_s1_write),                  //                                         .write
		.onchip_memory2_s1_readdata                     (mm_interconnect_0_onchip_memory2_s1_readdata),               //                                         .readdata
		.onchip_memory2_s1_writedata                    (mm_interconnect_0_onchip_memory2_s1_writedata),              //                                         .writedata
		.onchip_memory2_s1_byteenable                   (mm_interconnect_0_onchip_memory2_s1_byteenable),             //                                         .byteenable
		.onchip_memory2_s1_chipselect                   (mm_interconnect_0_onchip_memory2_s1_chipselect),             //                                         .chipselect
		.onchip_memory2_s1_clken                        (mm_interconnect_0_onchip_memory2_s1_clken),                  //                                         .clken
		.pio_height_s1_address                          (mm_interconnect_0_pio_height_s1_address),                    //                            pio_height_s1.address
		.pio_height_s1_readdata                         (mm_interconnect_0_pio_height_s1_readdata),                   //                                         .readdata
		.pio_key_s1_address                             (mm_interconnect_0_pio_key_s1_address),                       //                               pio_key_s1.address
		.pio_key_s1_write                               (mm_interconnect_0_pio_key_s1_write),                         //                                         .write
		.pio_key_s1_readdata                            (mm_interconnect_0_pio_key_s1_readdata),                      //                                         .readdata
		.pio_key_s1_writedata                           (mm_interconnect_0_pio_key_s1_writedata),                     //                                         .writedata
		.pio_key_s1_chipselect                          (mm_interconnect_0_pio_key_s1_chipselect),                    //                                         .chipselect
		.pio_led_s1_address                             (mm_interconnect_0_pio_led_s1_address),                       //                               pio_led_s1.address
		.pio_led_s1_write                               (mm_interconnect_0_pio_led_s1_write),                         //                                         .write
		.pio_led_s1_readdata                            (mm_interconnect_0_pio_led_s1_readdata),                      //                                         .readdata
		.pio_led_s1_writedata                           (mm_interconnect_0_pio_led_s1_writedata),                     //                                         .writedata
		.pio_led_s1_chipselect                          (mm_interconnect_0_pio_led_s1_chipselect),                    //                                         .chipselect
		.pio_width_s1_address                           (mm_interconnect_0_pio_width_s1_address),                     //                             pio_width_s1.address
		.pio_width_s1_readdata                          (mm_interconnect_0_pio_width_s1_readdata),                    //                                         .readdata
		.pio_wifi_reset_s1_address                      (mm_interconnect_0_pio_wifi_reset_s1_address),                //                        pio_wifi_reset_s1.address
		.pio_wifi_reset_s1_write                        (mm_interconnect_0_pio_wifi_reset_s1_write),                  //                                         .write
		.pio_wifi_reset_s1_readdata                     (mm_interconnect_0_pio_wifi_reset_s1_readdata),               //                                         .readdata
		.pio_wifi_reset_s1_writedata                    (mm_interconnect_0_pio_wifi_reset_s1_writedata),              //                                         .writedata
		.pio_wifi_reset_s1_chipselect                   (mm_interconnect_0_pio_wifi_reset_s1_chipselect),             //                                         .chipselect
		.pio_x_s1_address                               (mm_interconnect_0_pio_x_s1_address),                         //                                 pio_x_s1.address
		.pio_x_s1_readdata                              (mm_interconnect_0_pio_x_s1_readdata),                        //                                         .readdata
		.pio_y_s1_address                               (mm_interconnect_0_pio_y_s1_address),                         //                                 pio_y_s1.address
		.pio_y_s1_readdata                              (mm_interconnect_0_pio_y_s1_readdata),                        //                                         .readdata
		.SEG7_IF_0_avalon_slave_address                 (mm_interconnect_0_seg7_if_0_avalon_slave_address),           //                   SEG7_IF_0_avalon_slave.address
		.SEG7_IF_0_avalon_slave_write                   (mm_interconnect_0_seg7_if_0_avalon_slave_write),             //                                         .write
		.SEG7_IF_0_avalon_slave_read                    (mm_interconnect_0_seg7_if_0_avalon_slave_read),              //                                         .read
		.SEG7_IF_0_avalon_slave_readdata                (mm_interconnect_0_seg7_if_0_avalon_slave_readdata),          //                                         .readdata
		.SEG7_IF_0_avalon_slave_writedata               (mm_interconnect_0_seg7_if_0_avalon_slave_writedata),         //                                         .writedata
		.sysid_qsys_control_slave_address               (mm_interconnect_0_sysid_qsys_control_slave_address),         //                 sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata              (mm_interconnect_0_sysid_qsys_control_slave_readdata),        //                                         .readdata
		.timer_s1_address                               (mm_interconnect_0_timer_s1_address),                         //                                 timer_s1.address
		.timer_s1_write                                 (mm_interconnect_0_timer_s1_write),                           //                                         .write
		.timer_s1_readdata                              (mm_interconnect_0_timer_s1_readdata),                        //                                         .readdata
		.timer_s1_writedata                             (mm_interconnect_0_timer_s1_writedata),                       //                                         .writedata
		.timer_s1_chipselect                            (mm_interconnect_0_timer_s1_chipselect),                      //                                         .chipselect
		.wifi_uart0_s1_address                          (mm_interconnect_0_wifi_uart0_s1_address),                    //                            wifi_uart0_s1.address
		.wifi_uart0_s1_write                            (mm_interconnect_0_wifi_uart0_s1_write),                      //                                         .write
		.wifi_uart0_s1_read                             (mm_interconnect_0_wifi_uart0_s1_read),                       //                                         .read
		.wifi_uart0_s1_readdata                         (mm_interconnect_0_wifi_uart0_s1_readdata),                   //                                         .readdata
		.wifi_uart0_s1_writedata                        (mm_interconnect_0_wifi_uart0_s1_writedata),                  //                                         .writedata
		.wifi_uart0_s1_begintransfer                    (mm_interconnect_0_wifi_uart0_s1_begintransfer),              //                                         .begintransfer
		.wifi_uart0_s1_chipselect                       (mm_interconnect_0_wifi_uart0_s1_chipselect)                  //                                         .chipselect
	);

	RFS_WiFi_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
