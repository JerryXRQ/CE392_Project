module  painting_top(

	//////////// CLOCK //////////
	input 		          		FPGA_CLK1_50,
	input 		          		FPGA_CLK2_50,
	input 		          		FPGA_CLK3_50,	
	//////////// HDMI //////////
	inout 		          		HDMI_I2C_SCL,
	inout 		          		HDMI_I2C_SDA,
	inout 		          		HDMI_I2S,
	inout 		          		HDMI_LRCLK,
	inout 		          		HDMI_MCLK,
	inout 		          		HDMI_SCLK,
	output		          		HDMI_TX_CLK,
	output		          		HDMI_TX_DE,
	output		    [23:0]		HDMI_TX_D,
	output		          		HDMI_TX_HS,
	input 		          		HDMI_TX_INT,
	output		          		HDMI_TX_VS,

	//////////// KEY //////////
	input 		     [1:0]		KEY,

	//////////// LED //////////
	// output		     [7:0]		LED,

	//////////// SW //////////
	input 		     [3:0]		SW,

	//////////// GPIO_0, GPIO connect to D8M-GPIO //////////
	inout 		          		CAMERA_I2C_SCL,
	inout 		          		CAMERA_I2C_SDA,
	output		          		CAMERA_PWDN_n,
	output		          		MIPI_CS_n,
	inout 		          		MIPI_I2C_SCL,
	inout 		          		MIPI_I2C_SDA,
	output		          		MIPI_MCLK,
	input 		          		MIPI_PIXEL_CLK,
	input 		     [9:0]		MIPI_PIXEL_D,
	input 		          		MIPI_PIXEL_HS,
	input 		          		MIPI_PIXEL_VS,
	output		          		MIPI_REFCLK,
	output		          		MIPI_RESET_n
);

logic                       valid_out;

logic [7:0]		LED;


//assign FPGA_CLK1_50 = SYS_CLK;
//assign FPGA_CLK2_50 = SYS_CLK;
//assign FPGA_CLK3_50 = SYS_CLK;

//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

DE10_NANO_D8M_RTL DE10_NANO_D8M_RTL_INST(

	//////////// CLOCK //////////
	.FPGA_CLK1_50(FPGA_CLK1_50),
	.FPGA_CLK2_50(FPGA_CLK2_50),
	.FPGA_CLK3_50(FPGA_CLK3_50),

	//////////// HDMI //////////
	.HDMI_I2C_SCL(HDMI_I2C_SCL),
	.HDMI_I2C_SDA(HDMI_I2C_SDA),
	.HDMI_I2S(HDMI_I2S),
	.HDMI_LRCLK(HDMI_LRCLK),
	.HDMI_MCLK(HDMI_MCLK),
	.HDMI_SCLK(HDMI_SCLK),
	.HDMI_TX_CLK(HDMI_TX_CLK),
	.HDMI_TX_DE(HDMI_TX_DE),
	.HDMI_TX_D(HDMI_TX_D),
	.HDMI_TX_HS(HDMI_TX_HS),
	.HDMI_TX_INT(HDMI_TX_INT),
	.HDMI_TX_VS(HDMI_TX_VS),

	//////////// KEY //////////
	.KEY(KEY),

	//////////// LED //////////
	.LED(LED),

	//////////// SW //////////
	.SW(SW),

	//////////// GPIO_0, GPIO connect to D8M-GPIO //////////
	.CAMERA_I2C_SCL(CAMERA_I2C_SCL),
	.CAMERA_I2C_SDA(CAMERA_I2C_SDA),
	.CAMERA_PWDN_n(CAMERA_PWDN_n),
	.MIPI_CS_n(MIPI_CS_n),
	.MIPI_I2C_SCL(MIPI_I2C_SCL),
	.MIPI_I2C_SDA(MIPI_I2C_SDA),
	.MIPI_MCLK(MIPI_MCLK),
	.MIPI_PIXEL_CLK(MIPI_PIXEL_CLK),
	.MIPI_PIXEL_D(MIPI_PIXEL_D),
	.MIPI_PIXEL_HS(MIPI_PIXEL_HS),
	.MIPI_PIXEL_VS(MIPI_PIXEL_VS),
	.MIPI_REFCLK(MIPI_REFCLK),
	.MIPI_RESET_n(MIPI_RESET_n),

	//////////// tracking location //////////
	.valid_out(valid_out)
    // output			[11:0]		center_x_out,
    // output			[11:0]		center_y_out,
    // output			[11:0]		width_out,
    // output			[11:0]		height_out

);


//empty_test empty_test_inst(
//    .valid_out(valid_out)
//);

endmodule