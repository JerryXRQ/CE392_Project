
module empty_test (
    input  logic valid_out
);


endmodule